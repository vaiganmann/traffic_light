`include "counter.sv"

//the high level module
module traffic_light (output bit red_o, yellow_o, green_o,
             input bit clk_i, rst_i
             );

parameter period_red = 3, period_yellow_red = 3, period_yellow = 3, period_blinky_green = 3, period_green = 3;//number of cloks of a light
bit [10:0] nr = period_red, nyr = period_yellow_red, ny = period_yellow, nbg = period_blinky_green, ng = period_green;
bit [10:0] next_current_count, current_count, count ;
bit start, rst, overflow, current_green, next_current_green;
//****************************************************************
//            Some local defs
//****************************************************************
typedef enum {RST, RED,YELLOW_RED, GREEN, BLINKY_GREEN, YELLOW} states;
states next_state_t , state_t; 

counter counter_inst(clk_i, rst_i, count, current_count , overflow);

//****************************************************************
//            Finite State machine 
//****************************************************************
always_ff @(posedge clk_i or posedge rst_i) begin
    if (rst_i) begin
       state_t <= RST;
       current_count <= nr-1;
       current_green <= 0;
    end
      else begin
        state_t <= next_state_t;
        current_count <= next_current_count;
        current_green <= next_current_green;
      end
end

always_comb begin : set_next_state 
 
next_state_t = state_t;
next_current_count = current_count;

     unique case(state_t)
      RST: begin
            next_state_t = RED; 
            next_current_count = nr-1;
           end
      RED: begin      
            if (overflow)
              begin
                next_current_count = nyr-1;
                next_state_t = YELLOW_RED;
              end
            end        
      YELLOW_RED: begin              
              if (overflow)
                 begin
                    next_current_count = ng-1;
                    next_state_t = GREEN;
                 end
               end
      GREEN: begin             
              if (overflow)
                begin
				          next_current_count = nbg-1;
				          next_state_t = BLINKY_GREEN; 
                end
              end
      BLINKY_GREEN: begin
               if (overflow) 
                  begin
                    next_state_t =  YELLOW;
				            next_current_count = ny-1;
                end
               end
      YELLOW: begin
                if (overflow) begin
				          next_current_count = nr-1;
				          next_state_t =  RED;
                end
              end 
    endcase 
end:set_next_state

always_comb begin:set_outputs
next_current_green = current_green;
 {red_o, green_o, yellow_o} = 3'b000;
     unique case(state_t)
      RED:
        begin      
           red_o = 1;
        end      
      YELLOW_RED:
        begin              
            red_o = 1;
            yellow_o = 1;
        end
      GREEN: 
        begin
             green_o = 1;
        end
      BLINKY_GREEN: 
        begin
            if(!current_green)
                begin
                 green_o = 1;
                 next_current_green = 1;
                end
            else
              begin
                green_o = 0;
                next_current_green = 0;
              end
        end      
      YELLOW:
       begin
             yellow_o = 1;
       end 
    endcase 
end:set_outputs
endmodule 


module testbench;
bit clk_i, rst_i; 
bit red_o, yellow_o, green_o;  

 traffic_light #(.period_red(20)) DUT(.* , .rst_i(1'b0));

 
initial begin clk_i = 1'b0;
forever #10  clk_i = !clk_i;
end

endmodule

